
package mem_pkg;
  parameter int MEM_DEPTH = 1024;   // 1024 memory locations
  parameter int FIFO_DEPTH = 16;   // FIFO can hold 16 transactions

  //`include "axi_if.sv"
  //`include "axi_memory.sv"
endpackage
